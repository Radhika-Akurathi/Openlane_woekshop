*Model Description
.param temp=27


*Including sky130 library files
.lib "sky130_fd_pr/models/sky130.lib.spice" tt


*Netlist Description



XM1 Vdd n1 0 0 sky130_fd_pr__nfet_01v8 w=0.65 l=0.25

R1 in n1 55

Vdd vdd 0 1.8V
Vin in 0 1.8V

*simulation commands

.op 
.dc Vdd 0 1.8 0.1 Vin 0 1.8 0.2



.end

